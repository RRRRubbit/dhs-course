LIBRARY IEEE;
USE IEEE.ELECTRICAL_SYSTEMS.ALL;

ENTITY diode_E IS
  
  PORT (
    TERMINAL anode, cathode : ELECTRICAL);

END diode_E;

-- Architecture to be added by the students
